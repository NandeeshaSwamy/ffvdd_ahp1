`include "design.sv"
`include "transaction.sv"
`include "generator.sv"
`include "interface.sv"
`include "driver.sv"
`include "environment.sv"


`include "random_test.sv"


`include "testbench.sv"




