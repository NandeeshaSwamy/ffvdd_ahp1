
interface intf(input logic clk);
  
  //declaring the signals
  logic in;
  logic d0;
  logic d1;
  logic q0;
  logic q1;
  
endinterface
